library ieee ;
use ieee.std_logic_1164.all ;
entity reg6 is
   port ( resetN , clk : in  std_logic                      ;
          ena          : in  std_logic                      ;
          din          : in  std_logic_vector(5 downto 0)   ;
          dout         : out std_logic_vector(5 downto 0) ) ;
end reg6 ;
architecture arc_reg6 of reg6 is
begin
   process( resetN , clk )
   begin
      if resetN = '0' then
         dout <= "110000" ;
      elsif clk'event and clk = '1' then
         if ena = '1' then
            dout <= din ;
         end if ;
      end if ;
   end process ;
end arc_reg6 ;
   